module debouncer(
  input [3:0] digit, 
  output [6:0] cathode
)